module FP_divider_newfpu(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
`endif // RANDOMIZE_REG_INIT
  wire  FP_reciprocal_newfpu_clock; // @[FloatingPointDesigns.scala 2175:28]
  wire  FP_reciprocal_newfpu_reset; // @[FloatingPointDesigns.scala 2175:28]
  wire [31:0] FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2175:28]
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2178:28]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2178:28]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2178:28]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2178:28]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2178:28]
  reg [31:0] regs_0; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_1; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_2; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_3; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_4; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_5; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_6; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_7; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_8; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_9; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_10; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_11; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_12; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_13; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_14; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_15; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_16; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_17; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_18; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_19; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_20; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_21; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_22; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_23; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_24; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_25; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_26; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_27; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_28; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_29; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_30; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_31; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_32; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_33; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_34; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_35; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_36; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_37; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_38; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_39; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_40; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_41; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_42; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_43; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_44; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_45; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_46; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_47; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_48; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_49; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_50; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_51; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_52; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_53; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_54; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_55; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_56; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_57; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_58; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_59; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_60; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_61; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_62; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_63; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_64; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_65; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_66; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_67; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_68; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_69; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_70; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_71; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_72; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_73; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_74; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_75; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_76; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_77; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_78; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_79; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_80; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_81; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_82; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_83; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_84; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_85; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_86; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_87; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_88; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_89; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_90; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_91; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_92; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_93; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_94; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_95; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_96; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_97; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_98; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_99; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_100; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_101; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_102; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_103; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_104; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_105; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_106; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_107; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_108; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_109; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_110; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_111; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_112; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_113; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_114; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_115; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_116; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_117; // @[FloatingPointDesigns.scala 2170:23]
  reg [31:0] regs_118; // @[FloatingPointDesigns.scala 2170:23]
  FP_reciprocal_newfpu FP_reciprocal_newfpu ( // @[FloatingPointDesigns.scala 2175:28]
    .clock(FP_reciprocal_newfpu_clock),
    .reset(FP_reciprocal_newfpu_reset),
    .io_out_s(FP_reciprocal_newfpu_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2178:28]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  assign io_out_s = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2182:14]
  assign FP_reciprocal_newfpu_clock = clock;
  assign FP_reciprocal_newfpu_reset = reset;
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = regs_118; // @[FloatingPointDesigns.scala 2180:21]
  assign FP_multiplier_10ccs_io_in_b = FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2181:21]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_0 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_0 <= io_in_a; // @[FloatingPointDesigns.scala 2171:13]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_1 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_1 <= regs_0; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_2 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_2 <= regs_1; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_3 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_3 <= regs_2; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_4 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_4 <= regs_3; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_5 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_5 <= regs_4; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_6 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_6 <= regs_5; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_7 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_7 <= regs_6; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_8 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_8 <= regs_7; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_9 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_9 <= regs_8; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_10 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_10 <= regs_9; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_11 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_11 <= regs_10; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_12 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_12 <= regs_11; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_13 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_13 <= regs_12; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_14 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_14 <= regs_13; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_15 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_15 <= regs_14; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_16 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_16 <= regs_15; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_17 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_17 <= regs_16; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_18 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_18 <= regs_17; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_19 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_19 <= regs_18; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_20 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_20 <= regs_19; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_21 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_21 <= regs_20; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_22 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_22 <= regs_21; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_23 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_23 <= regs_22; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_24 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_24 <= regs_23; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_25 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_25 <= regs_24; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_26 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_26 <= regs_25; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_27 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_27 <= regs_26; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_28 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_28 <= regs_27; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_29 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_29 <= regs_28; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_30 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_30 <= regs_29; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_31 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_31 <= regs_30; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_32 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_32 <= regs_31; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_33 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_33 <= regs_32; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_34 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_34 <= regs_33; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_35 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_35 <= regs_34; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_36 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_36 <= regs_35; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_37 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_37 <= regs_36; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_38 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_38 <= regs_37; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_39 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_39 <= regs_38; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_40 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_40 <= regs_39; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_41 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_41 <= regs_40; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_42 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_42 <= regs_41; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_43 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_43 <= regs_42; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_44 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_44 <= regs_43; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_45 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_45 <= regs_44; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_46 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_46 <= regs_45; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_47 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_47 <= regs_46; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_48 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_48 <= regs_47; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_49 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_49 <= regs_48; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_50 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_50 <= regs_49; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_51 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_51 <= regs_50; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_52 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_52 <= regs_51; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_53 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_53 <= regs_52; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_54 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_54 <= regs_53; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_55 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_55 <= regs_54; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_56 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_56 <= regs_55; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_57 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_57 <= regs_56; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_58 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_58 <= regs_57; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_59 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_59 <= regs_58; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_60 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_60 <= regs_59; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_61 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_61 <= regs_60; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_62 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_62 <= regs_61; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_63 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_63 <= regs_62; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_64 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_64 <= regs_63; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_65 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_65 <= regs_64; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_66 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_66 <= regs_65; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_67 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_67 <= regs_66; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_68 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_68 <= regs_67; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_69 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_69 <= regs_68; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_70 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_70 <= regs_69; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_71 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_71 <= regs_70; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_72 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_72 <= regs_71; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_73 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_73 <= regs_72; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_74 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_74 <= regs_73; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_75 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_75 <= regs_74; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_76 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_76 <= regs_75; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_77 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_77 <= regs_76; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_78 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_78 <= regs_77; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_79 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_79 <= regs_78; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_80 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_80 <= regs_79; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_81 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_81 <= regs_80; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_82 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_82 <= regs_81; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_83 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_83 <= regs_82; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_84 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_84 <= regs_83; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_85 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_85 <= regs_84; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_86 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_86 <= regs_85; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_87 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_87 <= regs_86; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_88 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_88 <= regs_87; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_89 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_89 <= regs_88; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_90 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_90 <= regs_89; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_91 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_91 <= regs_90; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_92 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_92 <= regs_91; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_93 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_93 <= regs_92; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_94 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_94 <= regs_93; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_95 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_95 <= regs_94; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_96 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_96 <= regs_95; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_97 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_97 <= regs_96; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_98 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_98 <= regs_97; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_99 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_99 <= regs_98; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_100 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_100 <= regs_99; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_101 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_101 <= regs_100; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_102 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_102 <= regs_101; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_103 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_103 <= regs_102; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_104 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_104 <= regs_103; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_105 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_105 <= regs_104; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_106 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_106 <= regs_105; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_107 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_107 <= regs_106; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_108 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_108 <= regs_107; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_109 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_109 <= regs_108; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_110 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_110 <= regs_109; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_111 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_111 <= regs_110; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_112 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_112 <= regs_111; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_113 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_113 <= regs_112; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_114 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_114 <= regs_113; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_115 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_115 <= regs_114; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_116 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_116 <= regs_115; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_117 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_117 <= regs_116; // @[FloatingPointDesigns.scala 2173:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2170:23]
      regs_118 <= 32'h0; // @[FloatingPointDesigns.scala 2170:23]
    end else begin
      regs_118 <= regs_117; // @[FloatingPointDesigns.scala 2173:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  regs_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  regs_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  regs_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  regs_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  regs_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  regs_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  regs_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  regs_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  regs_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  regs_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  regs_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  regs_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  regs_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  regs_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  regs_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  regs_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  regs_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  regs_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  regs_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  regs_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  regs_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  regs_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  regs_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  regs_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  regs_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  regs_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  regs_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  regs_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  regs_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  regs_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  regs_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  regs_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  regs_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  regs_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  regs_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  regs_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  regs_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  regs_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  regs_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  regs_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  regs_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  regs_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  regs_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  regs_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  regs_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  regs_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  regs_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  regs_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  regs_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  regs_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  regs_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  regs_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  regs_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  regs_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  regs_118 = _RAND_118[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
